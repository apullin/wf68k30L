// ========================================================================
// Operand routing submodule
// ========================================================================
// ALU operand multiplexers, register file input muxes, bit field
// offset/width/BITPOS, branch prediction, and DBcc condition are all
// handled by the operand mux submodule.

    WF68K30L_OPERAND_MUX I_OPERAND_MUX (
        .CLK                    (CLK),
        .OP                     (OP),
        .OP_WB                  (OP_WB),
        .OP_SIZE                (OP_SIZE),
        .BIW_0                  (BIW_0),
        .BIW_0_WB_73            (BIW_0_WB_73),
        .BIW_1                  (BIW_1),
        .BIW_2                  (BIW_2),
        .ADR_MODE               (ADR_MODE),
        .PHASE2                 (PHASE2_MAIN),
        .DATA_TO_CORE           (DATA_TO_CORE),
        .DR_OUT_1               (DR_OUT_1),
        .DR_OUT_2               (DR_OUT_2),
        .AR_OUT_1               (AR_OUT_1),
        .AR_OUT_2               (AR_OUT_2),
        .ADR_EFF                (ADR_EFF),
        .PC                     (PC),
        .PC_EW_OFFSET           (PC_EW_OFFSET),
        .STATUS_REG             (STATUS_REG),
        .VBR                    (VBR),
        .CACR                   (CACR),
        .CAAR                   (CAAR),
        .SFC                    (SFC),
        .DFC                    (DFC),
        .MMU_SRP                (MMU_SRP),
        .MMU_CRP                (MMU_CRP),
        .MMU_TC                 (MMU_TC),
        .MMU_TT0                (MMU_TT0),
        .MMU_TT1                (MMU_TT1),
        .MMU_MMUSR              (MMU_MMUSR),
        .ALU_RESULT             (ALU_RESULT),
        .STORE_IDATA_B1         (STORE_IDATA_B1),
        .STORE_IDATA_B2         (STORE_IDATA_B2),
        .EXT_WORD               (EXT_WORD),
        .BUSY_MAIN              (BUSY_MAIN),
        .ADR_OFFSET_EXH         (ADR_OFFSET_EXH),
        .ADR_OFFSET_MAIN        (ADR_OFFSET_MAIN),
        .BUSY_EXH               (BUSY_EXH),
        .ALU_BSY                (ALU_BSY),
        .AR_WR_1                (AR_WR_1),
        .DR_WR_1                (DR_WR_1),
        .DFC_WR                 (DFC_WR),
        .SFC_WR                 (SFC_WR),
        .ISP_WR                 (ISP_WR),
        .MSP_WR                 (MSP_WR),
        .USP_WR                 (USP_WR),
        .FETCH_MEM_ADR          (FETCH_MEM_ADR),
        .USE_DREG               (USE_DREG),
        .VBR_RD                 (VBR_RD),
        .CACR_RD                (CACR_RD),
        .CAAR_RD                (CAAR_RD),
        .SFC_RD                 (SFC_RD),
        .DFC_RD                 (DFC_RD),
        .ISP_RD                 (ISP_RD),
        .MSP_RD                 (MSP_RD),
        .USP_RD                 (USP_RD),
        .MMU_SRP_RD             (MMU_SRP_RD),
        .MMU_CRP_RD             (MMU_CRP_RD),
        .MMU_TC_RD              (MMU_TC_RD),
        .MMU_TT0_RD             (MMU_TT0_RD),
        .MMU_TT1_RD             (MMU_TT1_RD),
        .MMU_MMUSR_RD           (MMU_MMUSR_RD),
        .SR_WR_EXH              (SR_WR_EXH),
        .ADn                    (ADn),
        .MOVEP_PNTR             (MOVEP_PNTR),
        .ALU_OP1_IN             (ALU_OP1_IN),
        .ALU_OP2_IN             (ALU_OP2_IN),
        .ALU_OP3_IN             (ALU_OP3_IN),
        .AR_IN_1                (AR_IN_1),
        .AR_IN_2                (AR_IN_2),
        .DR_IN_1                (DR_IN_1),
        .DR_IN_2                (DR_IN_2),
        .BF_OFFSET              (BF_OFFSET),
        .BF_WIDTH               (BF_WIDTH),
        .BITPOS                 (BITPOS),
        .BRANCH_ATN             (BRANCH_ATN),
        .DBcc_COND              (DBcc_COND),
        .DATA_IMMEDIATE         (DATA_IMMEDIATE),
        .ADR_OFFSET             (ADR_OFFSET)
    );
