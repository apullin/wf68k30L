// Routing section aggregator.
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_operand_mux.svh"
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_core_signals.svh"
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_bus_cache.svh"
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_misc_status.svh"
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_mmu_translate.svh"
`include "wf68k30L_top_sections/routing/wf68k30L_top_routing_bus_outputs.svh"
