// ---- Internal signal declarations ----
// File roadmap:
// 1) Flat signal declarations (grouped by role).
// 2) Helper functions (MMU/cache decode, match, and table-walk helpers).
// 3) Sequential state blocks (cache/MMU/register tracking).
// 4) Combinational routing (bus requests, translation, FC/CI/CBREQ generation).
// 5) Submodule instantiations and top-level glue muxes.
//
// Core pipeline, register-file, ALU, and bus control signals.

logic        ADn;
logic [31:0] ADR_CPY_EXH;
logic [31:0] ADR_EFF;
logic [31:0] ADR_EFF_WB;
logic [31:0] ADR_L;
logic [31:0] ADR_LATCH;
logic [2:0]  ADR_MODE;
logic [2:0]  ADR_MODE_MAIN;
logic        ADR_IN_USE;
logic [31:0] ADR_OFFSET;
logic [31:0] ADR_OFFSET_EXH;
logic [5:0]  ADR_OFFSET_MAIN;
logic [31:0] ADR_P;
logic [31:0] ADR_BUS_REQ_PHYS;
logic [31:0] ADR_P_PHYS;
logic [31:0] ADR_P_PHYS_CALC;
logic [31:0] ADR_P_PHYS_LATCH;
logic        ADR_MARK_UNUSED_MAIN;
logic        ADR_MARK_USED;
logic        AERR;
logic        ALU_ACK;
logic        ALU_BSY;
logic        ALU_COND;
logic        ALU_INIT;
logic        ALU_LOAD_OP1;
logic        ALU_LOAD_OP2;
logic        ALU_LOAD_OP3;
logic [31:0] ALU_OP1_IN;
logic [31:0] ALU_OP2_IN;
logic [31:0] ALU_OP3_IN;
logic        ALU_REQ;
logic [63:0] ALU_RESULT;
logic [2:0]  AMODE_SEL;
logic        AR_DEC;
logic [31:0] AR_IN_1;
logic [31:0] AR_IN_2;
logic        AR_IN_USE;
logic        AR_INC;
logic        AR_MARK_USED;
logic [31:0] AR_OUT_1;
logic [31:0] AR_OUT_2;
logic [2:0]  AR_SEL_RD_1;
logic [2:0]  AR_SEL_RD_1_MAIN;
logic [2:0]  AR_SEL_RD_2;
logic [2:0]  AR_SEL_WR_1;
logic [2:0]  AR_SEL_WR_2;
logic        AR_WR_1;
logic        AR_WR_2;
logic        AVECn_BUSIF;
logic        BERR_MAIN;
logic [4:0]  BITPOS;
logic [15:0] BIW_0;
logic [7:3]  BIW_0_WB_73;
logic [15:0] BIW_1;
logic [15:0] BIW_2;
logic [31:0] BF_OFFSET;
logic [5:0]  BF_WIDTH;
logic        BKPT_CYCLE;
logic        BKPT_INSERT;
logic        BRANCH_ATN;
logic        BUS_BSY;
logic        BUSY_EXH;
logic        BUSY_MAIN;
logic        BUSY_OPD;
logic        CC_UPDT;
logic [31:0] CAAR;
logic        CAAR_RD;
logic        CAAR_WR;
logic [31:0] CACR;
logic        CACR_RD;
logic        CACR_WR;
logic        CPU_SPACE;
logic        CPU_SPACE_EXH;
logic [2:0]  DFC;
logic        DFC_RD;
logic        DFC_WR;

// MMU programmer-visible registers and ATC/shadow structures.
logic [63:0] MMU_SRP;
logic [63:0] MMU_CRP;
logic [31:0] MMU_TC;
logic [31:0] MMU_TT0;
logic [31:0] MMU_TT1;
logic [31:0] MMU_MMUSR;
logic        MMU_TC_RD;
logic        MMU_TC_WR;
logic        MMU_SRP_RD;
logic        MMU_SRP_WR;
logic        MMU_CRP_RD;
logic        MMU_CRP_WR;
logic        MMU_TT0_RD;
logic        MMU_TT0_WR;
logic        MMU_TT1_RD;
logic        MMU_TT1_WR;
logic        MMU_MMUSR_RD;
logic        MMU_MMUSR_WR;
logic        MMU_ATC_FLUSH;
logic [31:0] MMU_ATC_FLUSH_COUNT;
localparam int MMU_ATC_LINES = 8;
logic [MMU_ATC_LINES-1:0] MMU_ATC_V;
logic [MMU_ATC_LINES-1:0] MMU_ATC_B;
logic [MMU_ATC_LINES-1:0] MMU_ATC_W;
logic [MMU_ATC_LINES-1:0] MMU_ATC_M;
logic [2:0]  MMU_ATC_FC [0:MMU_ATC_LINES-1];
logic [31:0] MMU_ATC_TAG[0:MMU_ATC_LINES-1];
logic [31:0] MMU_ATC_PTAG[0:MMU_ATC_LINES-1];
logic [$clog2(MMU_ATC_LINES)-1:0] MMU_ATC_REPL_PTR;
localparam int MMU_DESC_SHADOW_LINES = 256;
logic [MMU_DESC_SHADOW_LINES-1:0] MMU_DESC_SHADOW_V;
logic [31:0] MMU_DESC_SHADOW_ADDR[0:MMU_DESC_SHADOW_LINES-1];
logic [31:0] MMU_DESC_SHADOW_DATA[0:MMU_DESC_SHADOW_LINES-1];
logic [$clog2(MMU_DESC_SHADOW_LINES)-1:0] MMU_DESC_SHADOW_REPL_PTR;
logic        MMU_DESC_SHADOW_PENDING;
logic [31:0] MMU_DESC_SHADOW_PENDING_ADDR;
logic        MMU_DESC_SHADOW_PENDING_WR;

// Remaining datapath, handshake, trap, and runtime-translation signals.
logic        DR_WR_1;
logic        DR_WR_2;
logic        DR_MARK_USED;
logic [31:0] DATA_FROM_CORE;
logic [31:0] DATA;
logic [31:0] DATA_IN_EXH;
logic [31:0] DATA_IMMEDIATE;
logic [31:0] DATA_EXH;
logic        DATA_RD;
logic        DATA_WR;
logic        DATA_RD_EXH;
logic        DATA_WR_EXH;
logic        DATA_RD_MAIN;
logic        DATA_WR_MAIN;
logic        DATA_RDY;
logic        DATA_RDY_BUSIF;
logic        DATA_RDY_CACHE;
logic        MMU_FAULT_DATA_ACK;
logic        MMU_FAULT_OPCODE_ACK;
logic [31:0] DATA_TO_CORE;
logic [31:0] DATA_TO_CORE_BUSIF;
logic [31:0] DATA_TO_CORE_CACHE;
logic        DATA_LAST_FROM_CACHE;
logic        DATA_VALID;
logic        DATA_VALID_BUSIF;
logic        DATA_VALID_CACHE;
logic [31:0] DISPLACEMENT;
logic [31:0] DISPLACEMENT_MAIN;
logic [7:0]  DISPLACEMENT_EXH;
logic [31:0] DATA_BUFFER;
logic        DBcc_COND;
logic [31:0] DR_IN_1;
logic [31:0] DR_IN_2;
logic [31:0] DR_OUT_2;
logic [31:0] DR_OUT_1;
logic [2:0]  DR_SEL_WR_1;
logic [2:0]  DR_SEL_WR_2;
logic [2:0]  DR_SEL_RD_1;
logic [2:0]  DR_SEL_RD_2;
logic        DR_IN_USE;
logic        EW_ACK;
logic        EW_REQ_MAIN;
logic        EX_TRACE;
logic        EXEC_RDY;
logic        EXH_REQ;
logic [15:0] EXT_WORD;
logic [31:0] FAULT_ADR;
logic        FB;
logic        FC;
logic        FETCH_MEM_ADR;
logic [2:0]  FC_I;
logic [2:0]  FC_BUS_REQ;
logic [2:0]  FC_LATCH;
logic        HILOn;
logic [31:0] INBUFFER;
logic        INT_TRIG;
logic [2:0]  IPL;
logic        ISP_DEC;
logic        ISP_RD;
logic        ISP_LOAD_EXH;
logic        ISP_WR_MAIN;
logic        ISP_WR;
logic [9:0]  IVECT_OFFS;
logic        IPEND_In;
logic [2:0]  IRQ_PEND;
logic        IPIPE_FILL;
logic        IPIPE_FLUSH;
logic        IPIPE_FLUSH_EXH;
logic        IPIPE_FLUSH_MAIN;
logic        RTE_PIPE_LOAD;
logic [15:0] RTE_PIPE_BIW_0;
logic [15:0] RTE_PIPE_BIW_1;
logic [15:0] RTE_PIPE_BIW_2;
logic        RTE_PIPE_C_FAULT;
logic        RTE_PIPE_B_FAULT;
logic [2:0]  IPIPE_OFFESET;
logic        LOOP_BSY;
logic        LOOP_SPLIT;
logic        LOOP_EXIT;
int          MOVEP_PNTR;
logic        MSP_RD;
logic        MSP_WR;
logic        OPCODE_RD;
logic        OPCODE_RDY;
logic        OPCODE_RDY_BUSIF;
logic        OPCODE_RDY_BUSIF_CORE;
logic        OPCODE_VALID;
logic        OPCODE_VALID_BUSIF;
logic [15:0] OPCODE_TO_CORE;
logic [15:0] OPCODE_TO_CORE_BUSIF;
OP_SIZETYPE  OP_SIZE;
OP_SIZETYPE  OP_SIZE_BUS;
OP_SIZETYPE  OP_SIZE_EXH;
OP_SIZETYPE  OP_SIZE_MAIN;
OP_SIZETYPE  OP_SIZE_WB; // Writeback.
logic        OPCODE_REQ;
logic        OPCODE_REQ_CORE;
logic        OPCODE_REQ_I;
logic        OW_VALID;
logic        OPD_ACK_MAIN;
OP_68K       OP;
OP_68K       OP_WB;
logic        OW_REQ_MAIN;
logic [31:0] OUTBUFFER;
logic [31:0] PC;
logic        PHASE2_MAIN;
logic        PC_ADD_DISPL;
logic [7:0]  PC_ADR_OFFSET;
logic [3:0]  PC_EW_OFFSET;
logic        PC_INC;
logic        PC_INC_EXH;
logic        PC_INC_EXH_I;
logic [31:0] PC_L;
logic        PC_LOAD;
logic        PC_LOAD_EXH;
logic        PC_LOAD_MAIN;
logic [7:0]  PC_OFFSET;
logic [7:0]  PC_OFFSET_OPD;
logic        PC_RESTORE_EXH;
logic        RB;
logic        RC;
logic        RD_REQ;
logic        RD_REQ_I;
logic        DATA_RD_BUS;
logic        DATA_RDY_BUSIF_CORE;
logic        RMC;
logic        REFILLn_EXH;
logic        RESTORE_ISP_PC;
logic        RESET_CPU;
logic        RESET_IN;
logic        RESET_STRB;
logic        CIOUT_ASSERT;
logic        CBREQ_ASSERT;
logic        CBREQ_REQ_NOW;
logic        CBREQ_REQ_LATCH;
logic        CBREQ_INST_REQ_NOW;
logic        CBREQ_DATA_REQ_NOW;
logic        OPCODE_REQ_CORE_MISS;
logic        SP_ADD_DISPL;
logic        SP_ADD_DISPL_EXH;
logic        SP_ADD_DISPL_MAIN;
logic        SBIT;
logic [8:0]  SSW_80;
logic [2:0]  SFC;
logic        SFC_RD;
logic        SFC_WR;
logic [15:0] SR_CPY;
logic        SR_RD;
logic        SR_INIT;
logic        SR_CLR_MBIT;
logic        SR_WR;
logic        SR_WR_EXH;
logic        SR_WR_MAIN;
logic [3:0]  STACK_FORMAT;
int          STACK_POS;
logic [15:0] STATUS_REG;
logic        STATUSn_MAIN;
logic        STATUSn_EXH;
logic        STORE_ADR_FORMAT;
logic        STORE_ABS_HI;
logic        STORE_ABS_LO;
logic        STORE_AEFF;
logic        STORE_D16;
logic        STORE_D32_LO;
logic        STORE_D32_HI;
logic        STORE_DISPL;
logic        STORE_MEM_ADR;
logic        STORE_OD_HI;
logic        STORE_OD_LO;
logic        STORE_IDATA_B1;
logic        STORE_IDATA_B2;
logic        TRAP_AERR;
logic        TRAP_ILLEGAL;
TRAPTYPE_OPC TRAP_CODE_OPC;
logic        TRAP_cc;
logic        TRAP_CHK;
logic        TRAP_DIVZERO;
logic        TRAP_V;
logic        TRAP_MMU_CFG;
// Coprocessor interface model (HW-003 phase 4/5, no external coprocessor present).
logic [2:0]  CPIF_STATE;
logic        CPIF_ACTIVE;
logic [2:0]  CPIF_LAST_CAT;
logic [2:0]  CPIF_LAST_CPID;
logic [4:0]  CPIF_LAST_CIR;
logic [15:0] CPIF_LAST_OPWORD;
logic        CPIF_LAST_READ;
logic        CPIF_LAST_WRITE;
logic        CPIF_LAST_RESPONDED;
logic [4:0]  CPIF_LAST_RESP_CIR;
logic [3:0]  CPIF_LAST_PHASE_LEN;
logic [3:0]  CPIF_PHASE_STEPS_LEFT;
logic [3:0]  CPIF_RESP_DELAY_LEFT;
logic [3:0]  CPIF_STEP_INDEX;
logic [4:0]  CPIF_STEP_CIR;
logic        CPIF_STEP_READ;
logic        CPIF_STEP_WRITE;
logic [4:0]  CPIF_RESP_CIR_EXPECT;
logic        CPIF_REQ_PULSE;
logic        CPIF_STEP_PULSE;
logic        CPIF_RESP_PULSE;
logic        CPIF_NORESP_PULSE;
logic        CPIF_TIMEOUT_PULSE;
logic        CPIF_BADRESP_PULSE;
logic [31:0] CPIF_REQ_COUNT;
logic [31:0] CPIF_STEP_COUNT;
logic [31:0] CPIF_RESP_COUNT;
logic [31:0] CPIF_NORESP_COUNT;
logic [31:0] CPIF_TIMEOUT_COUNT;
logic [31:0] CPIF_BADRESP_COUNT;
logic [31:0] CPIF_PRIV_BYPASS_COUNT;
logic [31:0] CPIF_LINEF_NOPROTO_COUNT;
logic        CPIF_MODEL_EXC_ENABLE;
logic        CPIF_MODEL_EXC_ON_NORESP;
logic [1:0]  CPIF_MODEL_EXC_KIND;   // 0=pre, 1=mid, 2=post
logic [7:0]  CPIF_MODEL_EXC_VECTOR;
logic        CPIF_MODEL_RESP_ENABLE;
logic [3:0]  CPIF_MODEL_RESP_DELAY;
logic [4:0]  CPIF_MODEL_RESP_CIR;
logic        CPIF_TRAP_PRE;
logic        CPIF_TRAP_MID;
logic        CPIF_TRAP_POST;
logic [7:0]  CPIF_TRAP_VECTOR;
logic [31:0] CPIF_PRE_EXC_COUNT;
logic [31:0] CPIF_MID_EXC_COUNT;
logic [31:0] CPIF_POST_EXC_COUNT;
logic [31:0] CPIF_PROTO_COUNT;
logic        MMU_RUNTIME_REQ;
logic        MMU_RUNTIME_FAULT;
logic        MMU_RUNTIME_STALL;
logic        MMU_RUNTIME_ATC_REFILL;
logic [2:0]  MMU_RUNTIME_ATC_FC;
logic [31:0] MMU_RUNTIME_ATC_TAG;
logic [31:0] MMU_RUNTIME_ATC_PTAG;
logic        MMU_RUNTIME_ATC_B;
logic        MMU_RUNTIME_ATC_W;
logic        MMU_RUNTIME_ATC_M;
logic        MMU_WALK_DELAY_ARMED;
logic        UNMARK;
logic        USE_APAIR;
logic        USE_DFC;
logic        USE_SFC;
logic        USE_DPAIR;
logic        USE_DREG;
logic        USP_RD;
logic        USP_WR;
logic [31:0] VBR;
logic        VBR_WR;
logic        VBR_RD;
logic        WR_REQ;
logic        WR_REQ_I;

// Cache model state: instruction/data lookup, fill, and burst tracking.
logic        ICACHE_HIT_NOW;
logic        ICACHE_RDY;
logic [15:0] ICACHE_OPCODE_WORD;
logic        ICACHE_FILL_PENDING;
logic [31:0] ICACHE_FILL_ADDR;
logic        ICACHE_FILL_CACHEABLE;
logic [2:0]  ICACHE_FILL_FC;
logic        ICACHE_BURST_TRACK_VALID;
logic [3:0]  ICACHE_BURST_TRACK_LINE;
logic [23:0] ICACHE_BURST_TRACK_TAG;
logic        ICACHE_BURST_FILL_VALID;
logic [3:0]  ICACHE_BURST_FILL_LINE;
logic [23:0] ICACHE_BURST_FILL_TAG;
logic [7:0]  ICACHE_BURST_FILL_PENDING;
logic [2:0]  ICACHE_BURST_FILL_FC;
logic [2:0]  ICACHE_BURST_FILL_NEXT_WORD;
logic [23:0] ICACHE_TAG [0:15];
logic [7:0]  ICACHE_VALID [0:15];
logic [15:0] ICACHE_DATA [0:15][0:7];
logic        DCACHE_HIT_NOW;
logic [31:0] DCACHE_HIT_DATA_NOW;
logic        DCACHE_HIT_PENDING;
logic [31:0] DCACHE_HIT_DATA_PENDING;
logic [23:0] DCACHE_TAG [0:15];
logic [31:0] DCACHE_DATA [0:15][0:3];
logic [3:0]  DCACHE_VALID [0:15];
logic        DCACHE_READ_FILL_PENDING;
logic [31:0] DCACHE_READ_FILL_ADDR;
OP_SIZETYPE  DCACHE_READ_FILL_SIZE;
logic        DCACHE_READ_FILL_CACHEABLE;
logic [2:0]  DCACHE_READ_FILL_FC;
logic        DCACHE_BURST_TRACK_VALID;
logic [3:0]  DCACHE_BURST_TRACK_LINE;
logic [23:0] DCACHE_BURST_TRACK_TAG;
logic        DCACHE_BURST_FILL_VALID;
logic [3:0]  DCACHE_BURST_FILL_LINE;
logic [23:0] DCACHE_BURST_FILL_TAG;
logic [3:0]  DCACHE_BURST_FILL_PENDING;
logic [2:0]  DCACHE_BURST_FILL_FC;
logic [1:0]  DCACHE_BURST_FILL_NEXT_ENTRY;
logic        DCACHE_WRITE_PENDING;
logic [31:0] DCACHE_WRITE_ADDR;
OP_SIZETYPE  DCACHE_WRITE_SIZE;
logic [31:0] DCACHE_WRITE_DATA;
logic        DCACHE_WRITE_CACHEABLE;
logic        BURST_PREFETCH_OP_REQ;
logic        BURST_PREFETCH_DATA_REQ;
logic [2:0]  BURST_PREFETCH_OP_WORD;
logic [1:0]  BURST_PREFETCH_DATA_ENTRY;
logic [31:0] BURST_PREFETCH_ADDR;
logic [2:0]  BURST_PREFETCH_FC;
logic        BUS_CYCLE_BURST;
logic        BUS_CYCLE_BURST_IS_OP;
