// Helper section aggregator.
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_datapath.svh"
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_mmu_base.svh"
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_mmu_ptest.svh"
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_mmu_runtime_walk.svh"
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_cache.svh"
`include "wf68k30L_top_sections/helpers/wf68k30L_top_helpers_coprocessor.svh"
